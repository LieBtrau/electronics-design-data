BF494 (PSpice format)
.MODEL Q_BF494_N_1 NPN( BF=143.5 BR=1 IS=2.11F RB=10 RC=0 
+      CJC=9.631P VJC=750M MJC=330M TR=10N CJE=182.3P 
+      VJE=750M MJE=330M TF=612.1P EG=1.11 VAF=100 
+      XTB=2M KF=0 AF=1 )
.END
